module Processor();


endmodule