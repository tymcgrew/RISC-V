module Control();


endmodule